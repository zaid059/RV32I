`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11/10/2023 10:07:26 PM
// Design Name: 
// Module Name: inst_mem
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module inst_mem(
 input logic[31:0] A,
 input logic[31:0]WD,
 input logic clk,
 output logic[31:0]RD,
 input logic [3:0] WM
);
  // Memory for instructions
  logic [31:0] instr_memory[0:1023];
 
initial begin
  $readmemh("imem.mem",instr_memory);
end
assign RD=instr_memory[A[31:2]];
endmodule
